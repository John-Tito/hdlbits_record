module my_dff8 (
    input        clk,
    input  [7:0] d  ,
    output [7:0] q
);
endmodule
