module Countslow (
    input        clk    ,
    input        slowena,
    input        reset  ,
    output [3:0] q
);
    reg [3:0] q_a;
    always @(posedge clk ) begin
        if(reset == 1'b1 || ((q_a >= 9) && (slowena==1'b1)))
            q_a <= 4'h0;
        else
            begin
                if (slowena==1'b1)
                    q_a <= q_a + 4'h1;
                else
                    q_a <= q_a  ;
            end
    end
    assign q = q_a;
endmodule
