module my_dff (
    input  clk,
    input  d  ,
    output q
);
endmodule
