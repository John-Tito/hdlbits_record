module mod_a (
    output out1,
    output out2,
    input  in1 ,
    input  in2 ,
    input  in3 ,
    input  in4
);
endmodule
